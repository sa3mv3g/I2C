 
 //`include "main.v"
 
 module testbench;
	
	reg scl;
	reg sda;
	reg tb_flag;
	
	wire [7:0] data;
	wire tb_sda;
	
	I2C _i2c(scl, tb_sda, data);
		
	initial begin
		$dumpfile("main.vcd");
		$dumpvars(0,testbench);
	end

	assign tb_sda = sda;
	
initial begin
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;

// now reading
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b1; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b1;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b0; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b1; sda = 1'b0;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b1; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
#1 scl = 1'b0; sda = 1'bz;
end
 
 
 endmodule 
 